module UART_RX(
    
);
    
endmodule