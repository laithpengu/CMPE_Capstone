module UART_RX() begin
    
end